library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TB_InstructionDecoder is
end TB_InstructionDecoder;

architecture Behavioral of TB_InstructionDecoder is
    component InstructionDecoder
    port()

begin


end Behavioral;
