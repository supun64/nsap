library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Slow_Clk is
    Port ( Clk : out STD_LOGIC);
end Slow_Clk;

architecture Behavioral of Slow_Clk is

begin


end Behavioral;
